/////////////////////////////////
// Filename    : xlr8_servo.v
// Author      : Matt Weber
// Description : A collection of servo channels (up to 32) and the
//                AVR IO registers needed to access them.
//               The servos aren't completely independant. They are backed
//                by 16 timers and directly alias (e.g. servo[0] and [16] always
//                have the same pulse width, although they can be separately
//                enabled/disabled).
//                3 Registers
//                  ControlRegister : 
//                        [7]   = enable channel (strobe write, read=enable for selected channel)
//                        [6]   = disable channel (strobe, always read as zero)
//                        [5]   = update channel pulse width (strobe, always read as zero)
//                        [4:0] = servo channel to enable/disable/update
//                  PulseWidthL :  [7:0]= lower 8 bits of servo pulse width in microseconds
//                  PulseWidthH :  [3:0]= upper 4 bits of servo pulse width in microseconds
//                   There is a PulseWidth register pair for each servo channel. 
//                    When written, the channel to access is given in ControlReg[4:0].
//                    On write it sets the pulse width that will be set when the control
//                      register is written with the update bit set
//                    Read just returns the last value written, regardless of ControlReg[4:0]
//                   To start a channel typically the PulseWidth registers would be written
//                    first, then the control register with the desired channel indicated and
//                    both the enable and update bits set
//               Future work. It should be possible to measure pulse widths with very little
//                 additional hardware. On the rising edge of of a pin to be measured, store
//                 the value of timercnt into chan_pw[pin]. Then on the falling edge of the
//                 pin do chan_pw[pin] = timercnt - chan_pw[pin] and adjust for wrapping.
//                 For the pin that is selected by ControlReg[4:0], the value of chan_pw[pin]
//                 is copied into the PulseWidthH/L registers, except that while chan_pw[pin]
//                 is holding the rising edge time (i.e. the pin is high) PulseWidthH[7] is
//                 also set and the software library can use this to determine that it needs to
//                 read the register again to get a valid result.       
//
//               UPDATED June 2019 by Mike Berry
//                 Added additional parameter to control servo speed by using
//                 the upper 4 bits of SVPWH register (for easy backward
//                 compatibility) to define a speed of 1-15, where 15 is
//                 fastest, and 1 is the slowest setting (0 means go as fast
//                 as the servo is able, so effectively ignore the speed
//                 setting).  From a library perspective, the write and
//                 writeMicroseconds functions will need an extra (optional)
//                 speed parameter.
//
// Copyright 2015, Superion Technology Group. All Rights Reserved
/////////////////////////////////

module xlr8_servo
 #(parameter NUM_SERVOS = 12,
   parameter SVCR_ADDR  = 6'h0, // servo control register
   parameter SVPWH_ADDR = 6'h0, // servo pulse width high
   parameter SVPWL_ADDR = 6'h0) // servo pulse width low
  (input logic clk,
  input logic                   en1mhz, // clock enable at 1MHz rate
  input logic                   rstn,
  // Register access for registers in first 64
  input [5:0]                   adr,
  input [7:0]                   dbus_in,
  output [7:0]                  dbus_out,
  input                         iore,
  input                         iowe,
  output wire                   io_out_en,
  // Register access for registers not in first 64
  input wire [7:0]              ramadr,
  input wire                    ramre,
  input wire                    ramwe,
  input wire                    dm_sel,
  // External inputs/outputs
  output logic [NUM_SERVOS-1:0] servos_en,
  output logic [NUM_SERVOS-1:0] servos_out,
  input  logic [4:0]            priv_index,
  input logic                   priv_wr_pw,
  input logic [15:0]            priv_pw
  );

  /////////////////////////////////
  // Local Parameters
  /////////////////////////////////
  localparam NUM_TIMERS = (NUM_SERVOS <= 16) ? NUM_SERVOS : 16;
  // Registers in I/O address range x0-x3F (memory addresses -x20-0x5F)
  //  use the adr/iore/iowe inputs. Registers in the extended address
  //  range (memory address 0x60 and above) use ramadr/ramre/ramwe
  localparam  SVCR_DM_LOC   = (SVCR_ADDR >= 16'h60) ? 1 : 0;
  localparam  SVPWH_DM_LOC   = (SVPWH_ADDR >= 16'h60) ? 1 : 0;
  localparam  SVPWL_DM_LOC   = (SVPWL_ADDR >= 16'h60) ? 1 : 0;

  localparam SVEN_BIT   = 7;
  localparam SVDIS_BIT  = 6;
  localparam SVUP_BIT   = 5;
  localparam SVCHAN_LSB = 0;    

  /////////////////////////////////
  // Signals
  /////////////////////////////////
  /*AUTOREG*/
  /*AUTOWIRE*/ 
  logic svcr_sel;
  logic svpwh_sel;
  logic svpwl_sel;
  logic svcr_we ;
  logic svpwh_we ;
  logic svpwl_we ;
  logic svcr_re ;
  logic svpwh_re ;
  logic svpwl_re ;
  logic [7:0] svcr_rdata;
  logic       SVEN;
  logic [4:0] SVCHAN;
  logic [3:0] SVSPD;
  logic [3:0] SVPWH;
  logic [7:0] SVPWL;
  logic [4:0] chan_in;
  logic [11:0] chan_pw [NUM_SERVOS-1:0]; // pulse width per channel from SW
  logic [11:0] chan_pw_out [NUM_SERVOS-1:0]; // pulse width per channel to servos
  logic [3:0] chan_sp [NUM_SERVOS-1:0]; // servo speed per channel
  logic       pw_update [NUM_SERVOS-1:0]; // flag to indicate a pw update is safe
  logic [5:0] pw_chg [NUM_SERVOS-1:0]; //  increment/decrement value related to speed
  logic [14:0]  timercnt; // Need to count to 20000us. That's 15 bits.

  /////////////////////////////////
  // Functions and Tasks
  /////////////////////////////////

  /////////////////////////////////
  // Main Code
  /////////////////////////////////

  assign svcr_sel = SVCR_DM_LOC ?  (dm_sel && ramadr == SVCR_ADDR ) : (adr[5:0] == SVCR_ADDR[5:0] ); 
  assign svpwh_sel = SVPWH_DM_LOC ?  (dm_sel && ramadr == SVPWH_ADDR ) : (adr[5:0] == SVPWH_ADDR[5:0] );
  assign svpwl_sel = SVPWL_DM_LOC ?  (dm_sel && ramadr == SVPWL_ADDR ) : (adr[5:0] == SVPWL_ADDR[5:0] );
  assign svcr_we = svcr_sel && (SVCR_DM_LOC ?  ramwe : iowe); 
  assign svpwh_we = svpwh_sel && (SVPWH_DM_LOC ?  ramwe : iowe);
  assign svpwl_we = svpwl_sel && (SVPWL_DM_LOC ?  ramwe : iowe); 
  assign svcr_re = svcr_sel && (SVCR_DM_LOC ?  ramre : iore); 
  assign svpwh_re = svpwh_sel && (SVPWH_DM_LOC ?  ramre : iore);
  assign svpwl_re = svpwl_sel && (SVPWL_DM_LOC ?  ramre : iore); 

  assign dbus_out =  ({8{svcr_sel}} & svcr_rdata) |
                     ({8{svpwh_sel}} & {SVSPD,SVPWH}) | 
                     ({8{svpwl_sel}} & SVPWL); 
  assign io_out_en = svcr_re || 
                     svpwh_re ||
                     svpwl_re; 

   // Control Registers
  assign chan_in = dbus_in[SVCHAN_LSB +: 5];
  always @(posedge clk or negedge rstn) begin
    if (!rstn)  begin
      SVEN   <= 1'b0;
      SVCHAN <= 5'h0;
      servos_en <= {NUM_SERVOS{1'b0}};
    end else if (svcr_we) begin
      SVCHAN<= chan_in;
      SVEN  <= dbus_in[SVEN_BIT]  || 
                          (servos_en[chan_in] && ~dbus_in[SVDIS_BIT]);;
      servos_en[chan_in] <= dbus_in[SVEN_BIT] || 
                          (servos_en[chan_in] && ~dbus_in[SVDIS_BIT]);
    end else begin
      SVEN <= servos_en[SVCHAN];
    end
  end // always @ (posedge clk or negedge rstn)
  always @(posedge clk) begin
    if (svcr_we) begin
      // Max pulse we'll do is 2.4ms which is 2400 counts at 1MHz. Need 12 bits.
      if (dbus_in[SVUP_BIT])
        begin
          chan_pw[chan_in] <= {SVPWH,SVPWL};
          chan_sp[chan_in] <= SVSPD;
        end
    end
    if (priv_wr_pw)
      begin
        chan_pw[priv_index] <= priv_pw[11:0];
      end
  end // always @ (posedge clk or negedge rstn)
  assign svcr_rdata = ({7'h0,SVEN}   << SVEN_BIT) |
                      ({3'h0,SVCHAN} << SVCHAN_LSB);
  always @(posedge clk or negedge rstn) begin
    if (!rstn)  begin
      SVPWH <= 4'h0;
      SVSPD <= 4'h0;
    end else if (svpwh_we) begin
      SVPWH  <= dbus_in[3:0];
      SVSPD  <= dbus_in[7:4];
    end 
  end
  always @(posedge clk or negedge rstn) begin
    if (!rstn)  begin
      SVPWL <= 8'h0;
    end else if (svpwl_we) begin
      SVPWL  <= dbus_in;
    end
  end

  // Run the counter at 1MHz (divby16) for 1us resolution
  always @(posedge clk or negedge rstn) begin
    if (!rstn) begin
      /*AUTORESET*/
      // Beginning of autoreset for uninitialized flops
      timercnt <= 15'h0;
      // End of automatics
    end else if (en1mhz && |servos_en) begin
      // it takes 20000 cycles of 1MHz to get 20ms
      timercnt <= (timercnt == 15'd19999) ? 15'd0 : (timercnt + 15'd1);
    end
  end // always @ (posedge clk or negedge rstn)
  // Save gates by using common timer for all channels
  // By modifying 2 of the top 3 bits of the count, we can
  //  easily get up to four channels non-overlapping. Getting
  //  more to be non-overlapping is probably not worth the
  //  extra logic it would require.
  genvar i;
  generate 
    for (i=0;i<NUM_SERVOS;i++) begin : gen_chan
      // the increment/decrement value is 4X the chan_sp coming in
      assign pw_chg[i] = chan_sp[i] << 2;
      always @(posedge clk or negedge rstn) begin
        if (!rstn) begin
          servos_out[i] <= 1'b0;
          chan_pw_out[i] <= 12'd1500; // start centered then move
          pw_update[i] <= 1'b0; // avoid any glitches at startup
        end else begin
          // every 20ms (corresponds to every update of the servo pulse width)
          // update the value sent to to servo, incrementing or decrementing
          // based on the chan_sp value.
          //
          // Assume a nominal range of 1000-2000us, and assume the slowest
          // we'd want to go is 5 seconds.  20ms updates means 50/second, so
          // in 5 seconds we'll see 250 updates.  For 1000us of change, each
          // increment/decrement will be 4us for slowest operation, and 15X
          // that (since we have settings of 1-15) would be 60us per update
          // (which translates to 1/3 second for full travel).
          if ((chan_sp[i] == 4'd0) && pw_update[i]) begin
            chan_pw_out[i] <= chan_pw[i]; // pass the value through if chan_sp is zero
          end else if (en1mhz && (timercnt == 15'd0)) begin
            if (chan_pw[i] >= (chan_pw_out[i] + pw_chg[i])) begin
              chan_pw_out[i] <= chan_pw_out[i] + pw_chg[i];
            end else if (chan_pw[i] <= (chan_pw_out[i] - pw_chg[i])) begin
              chan_pw_out[i] <= chan_pw_out[i] - pw_chg[i];
            end else begin
              chan_pw_out[i] <= chan_pw[i];
            end
          end
          // Create the pw_update signal; set at timercnt==0; reset when timercnt>=chan_pw_out.
          // The purpose of this is to allow changes to chan_pw_out (for speed 0) any time during
          // an active pulse, but not after an output has gone low (this avoids a second runt
          // pulse during a single 20ms cycle).  This probably could be timercnt>chan_pw_out, but
          // if we're that close to the end, we'll play it conservative and shut 'er down.
          if (timercnt == 15'd0) begin
            pw_update[i] <= 1'b1;
          end else if (timercnt >= chan_pw_out[i]) begin
            pw_update[i] <= 1'b0;
          end
          // Do full less-than check instead of just checking for equals at the ends to 
          //  avoid missing a change in cases where chan_pw changes
          servos_out[i] <= servos_en[i] && (timercnt[14:12] == {1'b0,i[1:0]}) && (timercnt[11:0] <= chan_pw_out[i]);
        end
      end // always @ (posedge clk or negedge rstn)
    end // block: gen_chan
  endgenerate
  
   /////////////////////////////////
   // Assertions
   /////////////////////////////////

`ifdef STGI_ASSERT_ON
  assert property (@(posedge clk) disable iff (~rstn) (timercnt<=20000))
               else $display("ERROR: xlr8_servo : counter out of range");
`endif

   /////////////////////////////////
   // Cover Points
   /////////////////////////////////

`ifdef SUP_COVER_ON
`endif

endmodule

